--Include the standard library headers
library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Entity declaration
entity company_rework_2024_top is
    port(
        CLK                : in std_logic;
        RESET              : in std_logic;
        
        IN_VALID           : in std_logic;
        IN_START_OF_PACKET : in std_logic;
        IN_END_OF_PACKET   : in std_logic;
        IN_DATA            : in std_logic_vector(63 downto 0);
        IN_EMPTY           : in std_logic_vector(2 downto 0);
        IN_ERROR           : in std_logic;
        
        IN_READY           : out std_logic;
        OUT_VALID          : out std_logic;
        OUT_DATA           : out std_logic_vector(255 downto 0);
        OUT_BYTE_MASK      : out std_logic_vector(31 downto 0)
    );
end company_rework_2024_top;

--Architecture declaration
architecture rtl of company_rework_2024_top is
    --Signal declaration
    signal state         : std_logic_vector(2 downto 0);
    signal data          : std_logic_vector(255 downto 0);
    signal byte_mask     : std_logic_vector(31 downto 0);
    signal ready         : std_logic;
    signal out_valid     : std_logic;
    signal out_data      : std_logic_vector(255 downto 0);
    signal out_byte_mask : std_logic_vector(31 downto 0);

    --Added comment on testmp2 branch
    
    --Process declaration
    begin

end architecture rtl;
```